`ifndef _parameters_h
    `define _parameters_h
    localparam PROGRAM_MEMORY_SIZE_WORDS = 100;

    localparam REGISTER_WRITE_BYTE_UNSIGNED = 3'b 100;
    localparam REGISTER_WRITE_BYTE_SIGNED = 3'b 101;
    localparam REGISTER_WRITE_WORD = 3'b 010;
`endif
