`ifndef _parameters_h
`define _parameters_h
localparam PROGRAM_MEMORY_SIZE = 100; 
`endif
