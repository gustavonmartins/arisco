`default_nettype none
`include "rtl/utilities.v"

module consecutive_instructions_tb ();

reg clk;
reg reset;

SoC mut (
    .clk (clk), .reset (reset)
);
initial begin
    clk=0;
end
always begin
    #5;clk=~clk;
end

initial
begin
    $info("Unit testing consecutive instructions");
    $dumpfile("consecutive_instructions_tb.vcd");
    $dumpvars(0,mut);
    $monitor("%2t,reset=%b,clk=%b,pc=%d,current instruction=%h, state=%d",$time,reset,clk,mut.cpu.pc,mut.cpu.instruction,mut.cpu.single_instr.fsm_state);

    //I-Type instructions
    $info("Testing I-Type instructions");
    reset=1;#1;
    mut.rom.program_memory[0]={12'd 120, 5'd 0, 3'b 000, 5'd 5, 7'b 0010011};//imm[11:0] rs1 000 rd 0010011 I addi
    mut.rom.program_memory[1]={12'd 200, 5'd 0, 3'b 000, 5'd 5, 7'b 0010011};//imm[11:0] rs1 000 rd 0010011 I addi
    mut.rom.program_memory[2]={12'd 2000, 5'd 5, 3'b 000, 5'd 5, 7'b 0010011};//imm[11:0] rs1 000 rd 0010011 I addi
    mut.rom.program_memory[3]={12'b 111111111111, 5'd 0, 3'b 111, 5'd5, 7'b 0010011};// imm[11:0] rs1 111 rd 0010011 I andi
    mut.rom.program_memory[4]={12'b 1010,5'd 0,3'b 110,5'd 5,7'b 0010011}; // imm[11:0] rs1 110 rd 0010011 I ori
    @(negedge clk) #1;
    
    `resetFSMAndReadInstruction; // Resets FSM and reads first instruction2

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'd 120,"ADDI: Register 5 should contain 120");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'd 200,"ADDI: Register 5 should contain 200");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'd 2200,"ADDI: Register 5 should contain 2200");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'b 0,"ANDI: Register 5 should contain all zeroes");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'b 1010,"ORI: Register 5 should end with 1010");

    //R-Type instructions
    $info("Testing R-Type instructions");
    reset=1;#1;
    mut.rom.program_memory[0]={12'd 2,      5'd 0,  3'b 000,                5'd 29, 7'b 0010011};   //imm[11:0] rs1 000     rd  0010011     I addi
    mut.rom.program_memory[1]={12'd 5,      5'd 0,  3'b 000,                5'd 31, 7'b 0010011};   //imm[11:0] rs1 000     rd  0010011     I addi
    mut.rom.program_memory[2]={7'b 0,       5'd 29, 5'd 31,     3'b 000,    5'd 4,  7'b 0110011};   //0000000   rs2 rs1 000 rd  0110011  R add
    mut.rom.program_memory[3]={7'b 0100000, 5'd 29, 5'd 31,     3'b 000,    5'd 5,  7'b 0110011};   //0100000   rs2 rs1 000 rd  0110011  R sub
    mut.rom.program_memory[4]={12'd 2047,   5'd 0,  3'b 000,                5'd 10, 7'b 0010011};   //imm[11:0] rs1 000     rd  0010011     I addi
    mut.rom.program_memory[5]={12'd 2047,   5'd 0,  3'b 000,                5'd 11, 7'b 0010011};   //imm[11:0] rs1 000     rd  0010011     I addi
    mut.rom.program_memory[6]={7'b 0100000, 5'd 10, 5'd 11,     3'b 000,    5'd 6,  7'b 0110011};   //0100000   rs2 rs1 000 rd  0110011  R sub
    mut.rom.program_memory[7]={12'd 0,      5'd 0,  3'b 000,                5'd 0,  7'b 0010011};   //imm[11:0] rs1 000     rd  0010011     I addi NOOP
    
    @(negedge clk); @(negedge clk) #1; 
    
    reset=0;@(negedge clk);@(negedge clk);

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[29], 32'd 2,"ADDI: Register 29 should contain 2");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[31], 32'd 5,"ADDI: Register 31 should contain 5");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[4], 32'd 7,"ADD: Register 4 should contain 7");

    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[5], 32'd 3,"SUB: Register 5 should contain 3 = 5-2 ($31 - $29)");
    
    `fullFSMInstructionCycle // Just finished instruction
    `fullFSMInstructionCycle // Just finished instruction
    `fullFSMInstructionCycle // Just finished instruction
    `assertCaseEqual(mut.cpu.single_instr.reg_mem.memory[6], 32'd 0,"SUB: Register 6 should contain 0 = 2047 - 2 ($10 - $11)");

    #20;
    $display("Simulation finished");
    $finish;
end
endmodule
