`ifndef _parameters_h
`define _parameters_h
localparam PROGRAM_MEMORY_SIZE_WORDS = 100;
localparam MEMORY_SIZE_BYTES = 8192;
`endif
